module npu_write_buffer_manager(
    input   logic                       clk_i,
    input   logic                       rst_n,
    //command signal
    output  logic                       conv_finish_o,//convolution finish
    //ram interface
    output  logic   [15:0]              write_cs_o,//write chip select
    output  logic   [15:0][10:0]        write_addr_o,//write address
    output  logic   [15:0][127:0]       write_data_in_o,//write data
    output  logic   [15:0]              write_enable_o,//write enable
    output  logic   [15:0][15:0]        write_byte_enable_o,//write byte enable
    //configuration
    input   logic   [10:0]              reg_MEM_OUT_offset_x,
    input   logic   [3:0]               reg_MEM_OUT_offset_y,
    input   logic   [7:0]               reg_CONV_MODE_mode,//convolution mode
    input   logic   [11:0]              reg_FM_OCH_ST_och_st,//output channel start
    input   logic   [11:0]              reg_FM_OCH_ED_och_ed,//output channel end
    input   logic                       reg_CONV_MODE_full_ch,//full channel
    input   logic                       reg_CONV_MODE_ch_st,//full channel
    //from top
    input   logic                       en_i,//enable signal for whole npu
    //row_col_num_manager
    input   logic   [10:0]              nl_col_num_i,//column number from non-linear module
    input   logic   [10:0]              nl_row_num_i,//row number from non-linear module
    //from rbm
    input   logic   [7:0]               rbm_frame_num_i,//row frame from read buffer manager
    //datapath port
    input   logic   [3:0][7:0][15:0]    fm_in_i ,//input feature map
    input   logic                       fm_in_irdy_i,//input ready
    output  logic                       fm_in_trdy_o,//transform ready
    input   logic                       fm_in_last_i,//last signal for each row frame
    input   logic   [7:0]               fm_in_row_valid_i,//row valid signal
    input   logic   [3:0]               fm_in_ch_valid_i,//channel valid signal
    input   logic                       datapath_finish_i,//datapath finish signal
    input   logic                       row_frame_p//the possible additional row frame generated by pooling operation
);
localparam BYPASS = 8'h0;
localparam CONV3x3 = 8'h1;
localparam CONV3x3RGBA = 8'h2;
localparam CONV3x3DW = 8'h3;
localparam CONV1x1 = 8'h4;
localparam ELEMENTWISE_ADD = 8'h5;
localparam ELEMENTWISE_MUL = 8'h6;

logic   [17:0]              dividend_for_offset;//dividend for calculation of out_offset_x and out_offset_y
logic   [10:0]              out_offset_x;
logic   [10:0]              out_offset_y;

logic   [11:0]              wbm_och;
logic                       offset_half_entry;//the offset half entry in the first group

logic   [8:0]               num_half_group;//the number of half groups

logic                       last_col;//last column signal
logic                       last_frame;//last row frame signal
logic                       last_half_group;//last half group signal

logic   [3:0]               mem_start_index;//memory start index
logic   [3:0]               mem_end_index;//memory end index

logic   [15:0]              mem_col_start_1;//memory column start
logic   [15:0]              mem_col_start_2;

logic   [3:0]               num_valid_row;//number of valid rows
logic   [3:0]               valid_signal_2_ch;//valid for each 2 channels

logic   [7:0][3:0][15:0]    fm_in ;
logic   [15:0][7:0][15:0]   write_data_in ;

logic                       write_enable_cs, write_enable_ns;//write enable

logic   [15:0][3:0]         write_4byte_enable ;// one bit represent 16 bytes (8 channel)

logic   [15:0]              st_idx_plus_os_y;//start index plus offset y
logic   [15:0]              ed_idx_plus_os_y;//end index plus pffset y

logic                       wrap_around;//memory start index < memory end index

logic   [10:0]              write_addr_1;//write address
logic   [10:0]              write_addr_2;


//delay
logic   [3:0]               valid_signal_2_ch_d1;
logic                       fm_in_last_d1;
//fsm and sequential logic
enum logic [1:0] {IDLE, RUNNING} CS, NS;
logic   [10:0]              col_cs, col_ns;//current column
logic   [7:0]               curr_row_frame_cs, curr_row_frame_ns;//current row frame
logic                       curr_half_group_abs_cs, curr_half_group_abs_ns;//current half group absolute index in the matrix
logic   [10:0]              curr_half_group_cs, curr_half_group_ns;//current half group
logic   [15:0]              start_offset_cs, start_offset_ns;//offset of start_index and end_index
logic   [15:0]              start_index_cs, start_index_ns;//start index
logic   [15:0]              end_index_cs, end_index_ns;//end index
logic   [15:0]              write_chip_select_cs ;//write chip select
logic   [15:0]              write_chip_select_ns ;
logic   [15:0][10:0]        write_addr_cs ;//write address
logic   [15:0][10:0]        write_addr_ns ;
logic                       conv_finish_cs, conv_finish_ns;//convolution finish signal

assign dividend_for_offset = reg_FM_OCH_ST_och_st[11:4] * nl_row_num_i + reg_MEM_OUT_offset_y;
assign out_offset_x = reg_MEM_OUT_offset_x + dividend_for_offset[17:4] * nl_col_num_i;
assign out_offset_y = dividend_for_offset[3:0];

assign wbm_och = reg_FM_OCH_ED_och_ed - reg_FM_OCH_ST_och_st + 1;
// assign offset_half_entry = reg_FM_OCH_ST_och_st[4];
assign offset_half_entry = reg_FM_OCH_ST_och_st[3];
assign num_half_group = (wbm_och[2:0] == 3'b0) ? wbm_och[11:3] : (wbm_och[11:3] + 1);
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        fm_in_last_d1 <= 1'b0;
    end else begin
        if (NS == RUNNING && reg_CONV_MODE_full_ch == 1)begin
            if(!fm_in_irdy_i) begin
                fm_in_last_d1 <= fm_in_last_d1;
            end else begin
                fm_in_last_d1 <= fm_in_last_i;
            end
        end else begin
            fm_in_last_d1 <= 1'b0;
        end
    end
end
assign last_col = fm_in_last_d1;
assign last_frame = (curr_row_frame_cs == rbm_frame_num_i + row_frame_p - 1);
assign last_half_group = (curr_half_group_cs == num_half_group - 1);

always_comb begin
    if(fm_in_row_valid_i[7]) begin num_valid_row = 8; end
    else if(fm_in_row_valid_i[6]) begin num_valid_row = 7; end
    else if(fm_in_row_valid_i[5]) begin num_valid_row = 6; end
    else if(fm_in_row_valid_i[4]) begin num_valid_row = 5; end
    else if(fm_in_row_valid_i[3]) begin num_valid_row = 4; end
    else if(fm_in_row_valid_i[2]) begin num_valid_row = 3; end
    else if(fm_in_row_valid_i[1]) begin num_valid_row = 2; end
    else if(fm_in_row_valid_i[0]) begin num_valid_row = 1; end
    else begin num_valid_row = 0; end
end
always_comb begin
    if(curr_half_group_abs_ns == 0) begin
        valid_signal_2_ch[0] = (fm_in_ch_valid_i[1:0] == 2'b11);
        valid_signal_2_ch[1] = (fm_in_ch_valid_i[3:2] == 2'b11);
        valid_signal_2_ch[2] = 1'b0;
        valid_signal_2_ch[3] = 1'b0;
    end else begin
        valid_signal_2_ch[0] = 1'b0;
        valid_signal_2_ch[1] = 1'b0;
        valid_signal_2_ch[2] = (fm_in_ch_valid_i[1:0] == 2'b11);
        valid_signal_2_ch[3] = (fm_in_ch_valid_i[3:2] == 2'b11);
    end
end
always_comb begin
    case (CS)
        IDLE: begin
            if(fm_in_irdy_i) begin
                case (reg_CONV_MODE_mode)
                    CONV1x1, CONV3x3, CONV3x3RGBA, BYPASS, CONV3x3DW, ELEMENTWISE_ADD, ELEMENTWISE_MUL: begin
                        NS = RUNNING;
                    end
                    default: begin NS = IDLE; end
                endcase
            end else begin
                NS = CS;
            end
        end
        RUNNING: begin
            if (en_i == 0 || conv_finish_o) begin
                NS = IDLE;
            end else begin
                if(last_col == 1'b1 && last_frame == 1'b1 && last_half_group == 1'b1) begin
                    NS = IDLE;
                end else begin
                    NS = CS;
                end
            end
        end
        default: begin NS = IDLE; end
    endcase
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        CS <= IDLE;
    end else begin
        CS <= NS;
    end
end
always_comb begin
    if(CS == IDLE && NS == RUNNING) begin
        col_ns = 11'b0;
    end else begin
        if(!fm_in_irdy_i) begin
            col_ns = col_cs;
        end else begin
            case(CS)
                RUNNING: begin
                    if(last_col == 1'b1) begin
                        col_ns = 11'b0;
                    end else begin
                        col_ns = col_cs + 1;
                    end
                end
                default: begin col_ns = col_cs; end
            endcase
        end
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        col_cs <= 11'b0;
    end else begin
        col_cs <= col_ns;
    end
end
always_comb begin
    if(CS == IDLE && NS == RUNNING) begin
        curr_row_frame_ns = 8'b0;
    end else begin
        if(!fm_in_irdy_i) begin
            curr_row_frame_ns = curr_row_frame_cs;
        end else begin
            case (CS)
                RUNNING: begin
                    if(last_col == 1'b1 && last_frame == 1'b1) begin
                        curr_row_frame_ns = 8'b0;
                    end else if(last_col == 1'b1) begin
                        curr_row_frame_ns = curr_row_frame_cs + 1;
                    end else begin
                        curr_row_frame_ns = curr_row_frame_cs;
                    end
                end
                default: begin curr_row_frame_ns = curr_row_frame_cs; end
            endcase
        end
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        curr_row_frame_cs <= 8'b0;
    end else begin
        curr_row_frame_cs <= curr_row_frame_ns;
    end
end
always_comb begin
    if(CS == IDLE && NS == RUNNING) begin
        curr_half_group_abs_ns = offset_half_entry;
    end else begin
        if(!fm_in_irdy_i) begin
            curr_half_group_abs_ns = curr_half_group_abs_cs;
        end else begin
            case (CS)
                RUNNING: begin
                    curr_half_group_abs_ns = curr_half_group_ns[0] + offset_half_entry;
                end
                default: begin curr_half_group_abs_ns = curr_half_group_abs_cs; end
            endcase
        end
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        curr_half_group_abs_cs <= 1'b0;
    end else begin
        curr_half_group_abs_cs <= curr_half_group_abs_ns;
    end
end

always_comb begin
    if(CS == IDLE && NS == RUNNING) begin
        curr_half_group_ns = 11'b0;
    end else begin
        if(!fm_in_irdy_i) begin
            curr_half_group_ns = curr_half_group_cs;
        end else begin
            case (CS)
                RUNNING: begin
                    if(last_col == 1'b1 && last_frame == 1'b1 && last_half_group == 1'b1) begin
                        curr_half_group_ns = 11'b0;
                    end else if(last_col == 1'b1 && last_frame == 1'b1) begin
                        curr_half_group_ns = curr_half_group_cs + 1;
                    end else begin
                        curr_half_group_ns = curr_half_group_cs;
                    end
                end
                default: begin
                    curr_half_group_ns = curr_half_group_cs;
                end
            endcase
        end
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        curr_half_group_cs <= 11'b0;
    end else begin
        curr_half_group_cs <= curr_half_group_ns;
    end
end

always_comb begin
    if(CS == IDLE && NS == RUNNING) begin
        start_offset_ns = 16'b0;
    end else begin
        if(!fm_in_irdy_i) begin
            start_offset_ns = start_offset_cs;
        end else begin
            case (CS)
                RUNNING: begin
                    if(last_col == 1'b1 && last_frame == 1'b1 && last_half_group == 1'b1) begin
                        start_offset_ns = 16'b0;
                    end else if(last_col == 1'b1 && last_frame == 1'b1 && curr_half_group_abs_cs == 1'b1) begin
                        start_offset_ns = end_index_cs + 1;
                    end else begin
                        start_offset_ns = start_offset_cs;
                    end
                end
                default: begin
                    start_offset_ns = start_offset_cs;
                end
            endcase
        end
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        start_offset_cs <= 16'b0;
    end else begin
        start_offset_cs <= start_offset_ns;
    end
end

always_comb begin
    if(CS == IDLE && NS == RUNNING) begin
        if(!fm_in_irdy_i) begin
            write_enable_ns = 1'b0;
        end else begin
            write_enable_ns = 1'b1;
        end
    end else begin
        if(fm_in_irdy_i == 0 || fm_in_ch_valid_i == 0 || fm_in_row_valid_i == 0) begin
            write_enable_ns = 1'b0;
        end else begin
            case (CS)
                RUNNING: begin write_enable_ns = 1'b1; end
                default: begin write_enable_ns = 1'b0; end
            endcase
        end
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        write_enable_cs <= 1'b0;
    end else begin
        write_enable_cs <= write_enable_ns;
    end
end
always_comb begin
    if(CS == IDLE && NS == RUNNING) begin
        start_index_ns = 16'b0;
    end else begin
        if(!fm_in_irdy_i) begin
            start_index_ns = start_index_cs;
        end else begin
            case (CS)
                RUNNING: begin
                    if(last_col == 1'b1) begin
                        if(last_frame == 1'b1) begin
                            start_index_ns = start_offset_ns;
                        end else begin
                            start_index_ns = end_index_cs + 1;
                        end
                    end else begin
                        start_index_ns = start_index_cs;
                    end
                end
                default: begin start_index_ns = start_index_cs; end
            endcase
        end
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        start_index_cs <= 16'b0;
    end else begin
        start_index_cs <= start_index_ns;
    end
end
always_comb begin
    if(!fm_in_irdy_i) begin
        end_index_ns = end_index_cs;
    end else begin
        case (NS)
            RUNNING: begin
                end_index_ns = start_index_ns + num_valid_row - 1;
            end
            default: begin
                end_index_ns = end_index_cs;
            end
        endcase
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        end_index_cs <= 16'b0;
    end else begin
        end_index_cs <= end_index_ns;
    end
end

assign st_idx_plus_os_y = start_index_cs + out_offset_y;
assign ed_idx_plus_os_y = end_index_cs + out_offset_y;

assign mem_start_index = st_idx_plus_os_y[3:0];
assign mem_end_index = ed_idx_plus_os_y[3:0];

assign mem_col_start_1 = st_idx_plus_os_y[15:4] * nl_col_num_i + out_offset_x;
assign mem_col_start_2 = ed_idx_plus_os_y[15:4] * nl_col_num_i + out_offset_x;

assign wrap_around = mem_start_index > mem_end_index;

assign write_addr_1 = mem_col_start_1 + col_cs;
assign write_addr_2 = mem_col_start_2 + col_cs;

always_comb begin
    for(int unsigned i=0;i<16;i++) begin
        if(write_enable_cs == 1'b1) begin
            if(wrap_around == 1'b1) begin
                if(i >= mem_start_index) begin
                    write_addr_ns[i] = write_addr_1;
                    write_chip_select_ns[i] = 1'b1;
                end else if(i <= mem_end_index) begin
                    write_addr_ns[i] = write_addr_2;
                    write_chip_select_ns[i] = 1'b1;
                end else begin
                    write_addr_ns[i] = write_addr_cs[i];
                    write_chip_select_ns[i] = 1'b0;
                end
            end else begin
                if(i >= mem_start_index && i <= mem_end_index) begin
                    write_addr_ns[i] = write_addr_1;
                    write_chip_select_ns[i] = 1'b1;
                end else begin
                    write_addr_ns[i] = write_addr_cs[i];
                    write_chip_select_ns[i] = 1'b0;
                end
            end
        end else begin
            write_addr_ns[i] = write_addr_cs[i];
            write_chip_select_ns[i] = 1'b0;
        end
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        for(int i=0;i<16;i++) begin
            write_addr_cs[i] <= 11'b0;
            write_chip_select_cs[i] <= 1'b0;
        end
    end else begin
        for(int i=0;i<16;i++) begin
            write_addr_cs[i] <= write_addr_ns[i];
            write_chip_select_cs[i] <= write_chip_select_ns[i];
        end
    end
end
always_comb begin
    for(int i=0;i<16;i++) begin
        write_addr_o[i] = write_addr_cs[i];
        write_cs_o[i] = write_chip_select_cs[i];
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        for(int i=0;i<8;i++) begin
            for(int j=0;j<4;j++) begin
                fm_in[i][j] <= 16'b0;
            end
        end
    end else begin
        for(int i=0;i<8;i++) begin
            for(int j=0;j<4;j++) begin
                if(write_enable_ns) begin
                //notice there is a reverse of i and j
                    fm_in[i][j] <= fm_in_i[j][i];
                end else begin
                    fm_in[i][j] <= fm_in[i][j];
                end
            end
        end
    end
end

always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        valid_signal_2_ch_d1 <= 4'b0;
    end else begin
        valid_signal_2_ch_d1 <= valid_signal_2_ch;
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        for(int i=0;i<16;i++) begin
            for(int j=0;j<8;j++) begin
                write_data_in[i][j] <= 16'b0;
            end
        end
    end else begin
        for(int i=0;i<16;i++) begin
            for(int j=0;j<8;j++) begin
                if(write_enable_cs) begin
                    if(i < 8 && j < 4) begin
                        case ({curr_half_group_abs_cs, mem_start_index})
                            5'h00: begin write_data_in[i%16][j]         <= fm_in[i][j]; end
                            5'h01: begin write_data_in[(i+1)%16][j]     <= fm_in[i][j]; end
                            5'h02: begin write_data_in[(i+2)%16][j]     <= fm_in[i][j]; end
                            5'h03: begin write_data_in[(i+3)%16][j]     <= fm_in[i][j]; end
                            5'h04: begin write_data_in[(i+4)%16][j]     <= fm_in[i][j]; end
                            5'h05: begin write_data_in[(i+5)%16][j]     <= fm_in[i][j]; end
                            5'h06: begin write_data_in[(i+6)%16][j]     <= fm_in[i][j]; end
                            5'h07: begin write_data_in[(i+7)%16][j]     <= fm_in[i][j]; end
                            5'h08: begin write_data_in[(i+8)%16][j]     <= fm_in[i][j]; end
                            5'h09: begin write_data_in[(i+9)%16][j]     <= fm_in[i][j]; end
                            5'h0a: begin write_data_in[(i+10)%16][j]    <= fm_in[i][j]; end
                            5'h0b: begin write_data_in[(i+11)%16][j]    <= fm_in[i][j]; end
                            5'h0c: begin write_data_in[(i+12)%16][j]    <= fm_in[i][j]; end
                            5'h0d: begin write_data_in[(i+13)%16][j]    <= fm_in[i][j]; end
                            5'h0e: begin write_data_in[(i+14)%16][j]    <= fm_in[i][j]; end
                            5'h0f: begin write_data_in[(i+15)%16][j]    <= fm_in[i][j]; end
                            5'h10: begin write_data_in[i%16][j+4]      <= fm_in[i][j]; end
                            5'h11: begin write_data_in[(i+1)%16][j+4]  <= fm_in[i][j]; end
                            5'h12: begin write_data_in[(i+2)%16][j+4]  <= fm_in[i][j]; end
                            5'h13: begin write_data_in[(i+3)%16][j+4]  <= fm_in[i][j]; end
                            5'h14: begin write_data_in[(i+4)%16][j+4]  <= fm_in[i][j]; end
                            5'h15: begin write_data_in[(i+5)%16][j+4]  <= fm_in[i][j]; end
                            5'h16: begin write_data_in[(i+6)%16][j+4]  <= fm_in[i][j]; end
                            5'h17: begin write_data_in[(i+7)%16][j+4]  <= fm_in[i][j]; end
                            5'h18: begin write_data_in[(i+8)%16][j+4]  <= fm_in[i][j]; end
                            5'h19: begin write_data_in[(i+9)%16][j+4]  <= fm_in[i][j]; end
                            5'h1a: begin write_data_in[(i+10)%16][j+4] <= fm_in[i][j]; end
                            5'h1b: begin write_data_in[(i+11)%16][j+4] <= fm_in[i][j]; end
                            5'h1c: begin write_data_in[(i+12)%16][j+4] <= fm_in[i][j]; end
                            5'h1d: begin write_data_in[(i+13)%16][j+4] <= fm_in[i][j]; end
                            5'h1e: begin write_data_in[(i+14)%16][j+4] <= fm_in[i][j]; end
                            5'h1f: begin write_data_in[(i+15)%16][j+4] <= fm_in[i][j]; end
                        endcase
                    end
                end else begin
                    write_data_in[i][j] <= write_data_in[i][j];
                end
            end
        end
    end
end

always_comb begin
    for(int i=0;i<16;i++) begin
        for(int j=0;j<8;j++) begin
            for(int k=0;k<16;k++) begin
                write_data_in_o [i][16*j+k] = write_data_in[i][j][k];
            end
        end
    end
end

always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        for(int i=0;i<16;i++) begin
            for(int j=0;j<4;j++) begin
                write_4byte_enable[i][j] <= 1'b0;
            end
        end
    end else begin
        for(int i=0;i<16;i++) begin
            for(int j=0;j<4;j++) begin
                if(write_chip_select_ns[i] == 1'b1) begin
                    write_4byte_enable[i][j] <= valid_signal_2_ch_d1[j];
                end else begin
                    write_4byte_enable[i][j] <= 1'b0;
                end
            end
        end
    end
end
always_comb begin
    for(int i=0;i<16;i++) begin
        for(int j=0;j<4;j++) begin
            for(int k=0;k<4;k++) begin
                write_byte_enable_o[i][4*j+k] = write_4byte_enable[i][j];
            end
        end
    end
end

assign write_enable_o = write_cs_o;

assign fm_in_trdy_o = 1'b1;

// always_comb begin
//     if(last_col == 1'b1 && last_frame == 1'b1 && last_half_group == 1'b1) begin
//         conv_finish_ns <= 1'b1;
//     end else begin
//         conv_finish_ns <= 1'b0;
//     end
// end
// always_ff @(negedge rst_n, posedge clk_i) begin
//     if(!rst_n) begin
//         conv_finish_cs <= 1'b0;
//     end else begin
//         conv_finish_cs <= conv_finish_ns;
//     end
// end
// always_comb begin
//     if(reg_CONV_MODE_full_ch == 1'b1) begin
//         conv_finish_o = conv_finish_cs;
//     end else begin
//         conv_finish_o = datapath_finish_i;
//     end
// end

logic conv_finish_flag;
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        conv_finish_flag <= 1'b0;
    end else begin
        if(reg_CONV_MODE_full_ch == 1'b1 && (datapath_finish_i ^ conv_finish_cs))begin
            conv_finish_flag <= ~conv_finish_flag;
        end else begin
            conv_finish_flag <= conv_finish_flag;
        end 
    end
end

always_comb begin
    if(last_col == 1'b1 && last_frame == 1'b1 && last_half_group == 1'b1) begin
        conv_finish_ns <= 1'b1;
    end else begin
        conv_finish_ns <= 1'b0;
    end
end
always_ff @(negedge rst_n, posedge clk_i) begin
    if(!rst_n) begin
        conv_finish_cs <= 1'b0;
    end else begin
        conv_finish_cs <= conv_finish_ns;
    end
end
always_comb begin
    if(reg_CONV_MODE_full_ch == 1'b1) begin
        conv_finish_o = conv_finish_cs;
    end else begin
        conv_finish_o = datapath_finish_i;
    end
end

endmodule